
module Napot_Addr_Decode_Tb;

    Napot_Addr_Decode Napot_Addr_Decode_Inst();



endmodule